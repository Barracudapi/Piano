`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/12/02 17:40:03
// Design Name: 
// Module Name: clock1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module clock2(
input wire clk,rst,
output reg clk_1
    );
    //this is a clock divider
    //which output a clk with 0.5s period
    `include "ppppparameters.v"
    reg [31:0] div_cnt;
    
    
    always @(posedge clk, negedge rst) begin
        if(~rst)
            div_cnt <= 0;
        else if(div_cnt == TIME_075SEC) 
            div_cnt <= 0;
        else 
            div_cnt <= div_cnt + 1;
    end

    always @(posedge clk, negedge rst) begin
        if(~rst)
            clk_1 <= 0;
        else if( div_cnt == (TIME_075SEC>>1) -1)
            clk_1 <= 1;
        else if(div_cnt == TIME_075SEC -1 ) 
            clk_1 <= 0;
    end
    
    
    

endmodule
